module hello_world_top;
  initial begin
    $display("MESSI RULES THE WORLD!!");
    $display("OTHER");
  end
endmodule
